//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "somma_di_quadrati.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] B;    //: /sn:0 {0}(#:357,97)(357,126){1}
//: {2}(#:355,128)(316,128)(316,63){3}
//: {4}(357,130)(357,150){5}
reg enable;    //: /sn:0 {0}(78,307)(115,307){1}
supply0 w3;    //: /sn:0 {0}(414,528)(414,510){1}
reg [3:0] A;    //: /sn:0 {0}(#:217,97)(217,126){1}
//: {2}(217,126)(217,123)(217,123)(217,150){3}
//: {4}(#:215,128)(177,128)(177,63){5}
reg Clock;    //: /sn:0 {0}(6,196)(28,196){1}
//: {2}(32,196)(183,196){3}
//: {4}(30,194)(30,25)(282,25)(282,196)(323,196){5}
//: {6}(30,198)(30,270){7}
//: {8}(32,272)(115,272){9}
//: {10}(30,274)(30,523)(254,523){11}
wire [8:0] w0;    //: /sn:0 {0}(416,434)(#:416,405){1}
wire [7:0] w12;    //: /sn:0 {0}(#:283,472)(283,459){1}
//: {2}(285,457)(349,457){3}
//: {4}(353,457)(381,457){5}
//: {6}(351,455)(351,414){7}
//: {8}(283,455)(#:283,441){9}
wire w8;    //: /sn:0 {0}(249,300)(200,300)(200,300)(185,300){1}
wire [3:0] w2;    //: /sn:0 {0}(#:216,218)(216,236){1}
//: {2}(218,238)(#:267,238)(267,264){3}
//: {4}(214,238)(175,238)(175,218)(148,218){5}
wire [7:0] w15;    //: /sn:0 {0}(#:319,488)(346,488){1}
//: {2}(350,488)(#:381,488){3}
//: {4}(348,490)(#:348,500)(348,500)(348,556){5}
wire [3:0] w5;    //: /sn:0 {0}(#:356,218)(356,235){1}
//: {2}(#:358,237)(571,237)(571,227){3}
//: {4}(354,237)(#:300,237)(300,264){5}
wire [3:0] w9;    //: /sn:0 {0}(#:303,380)(303,349)(286,349){1}
//: {2}(284,347)(284,330){3}
//: {4}(282,349)(#:265,349)(#:265,380){5}
//: {6}(284,347)(#:284,357)(467,357)(467,318){7}
//: enddecls

  REG8bit g4 (.in(w12), .clk(Clock), .out(w15));   //: @(255, 473) /sz:(63, 64) /sn:0 /p:[ Ti0>0 Li0>11 Ro0<0 ]
  //: LED A0 (A) @(177,56) /sn:0 /w:[ 5 ] /type:3
  //: joint g8 (B) @(357, 128) /w:[ -1 1 2 4 ]
  //: LED g16 (w2) @(141,218) /sn:0 /R:1 /w:[ 5 ] /type:3
  MUL4x4 g3 (.a(w9), .b(w9), .p(w12));   //: @(251, 381) /sz:(65, 59) /R:3 /sn:0 /p:[ Ti0>5 Ti1>0 Bo0<9 ]
  //: DIP B (B) @(357,87) /sn:0 /w:[ 0 ] /st:15 /dn:1
  //: SWITCH enable (enable) @(61,307) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: joint g17 (w2) @(216, 238) /w:[ 2 1 4 -1 ]
  MUX4bit g2 (.b(w5), .a(w2), .c(w8), .out(w9));   //: @(250, 265) /sz:(68, 64) /sn:0 /p:[ Ti0>5 Ti1>3 Li0>0 Bo0<3 ]
  REG4bit g1 (.in(B), .clk(Clock), .out(w5));   //: @(324, 151) /sz:(68, 66) /sn:0 /p:[ Ti0>5 Li0>5 Bo0<0 ]
  //: DIP A (A) @(217,87) /sn:0 /w:[ 0 ] /st:15 /dn:1
  //: LED g18 (w9) @(467,311) /sn:0 /w:[ 7 ] /type:3
  //: joint g10 (w12) @(283, 457) /w:[ 2 8 -1 1 ]
  //: SWITCH Clock (Clock) @(-11,196) /sn:0 /w:[ 0 ] /st:1 /dn:1
  myCU g6 (.enable(enable), .clk(Clock), .c(w8));   //: @(116, 253) /sz:(68, 75) /sn:0 /p:[ Li0>1 Li1>9 Ro0<1 ]
  //: joint g7 (A) @(217, 128) /w:[ 2 1 4 -1 ]
  //: joint g9 (w9) @(284, 349) /w:[ 1 2 4 6 ]
  //: joint g22 (w15) @(348, 488) /w:[ 2 -1 1 4 ]
  //: joint g12 (Clock) @(30, 272) /w:[ 8 7 -1 10 ]
  //: LED g14 (w5) @(571,220) /sn:0 /w:[ 3 ] /type:3
  RCA8bit g5 (.b(w12), .a(w15), .C0(w3), .out(w0));   //: @(382, 435) /sz:(67, 75) /sn:0 /p:[ Li0>5 Li1>3 Bi0>1 To0<0 ]
  //: GROUND g11 (w3) @(414,534) /sn:0 /w:[ 0 ]
  //: LED g21 (w15) @(348,563) /sn:0 /R:2 /w:[ 5 ] /type:3
  //: LED g19 (w12) @(351,407) /sn:0 /w:[ 7 ] /type:3
  //: joint g20 (w12) @(351, 457) /w:[ 4 6 3 -1 ]
  //: joint g15 (w5) @(356, 237) /w:[ 2 1 4 -1 ]
  REG4bit g0 (.in(A), .clk(Clock), .out(w2));   //: @(184, 151) /sz:(68, 66) /sn:0 /p:[ Ti0>3 Li0>3 Bo0<0 ]
  //: LED ris (w0) @(416,398) /sn:0 /w:[ 1 ] /type:3
  //: LED B0 (B) @(316,56) /sn:0 /w:[ 3 ] /type:3
  //: joint g13 (Clock) @(30, 196) /w:[ 2 4 1 6 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDls
module FFDls(q, clk, D);
//: interface  /sz:(61, 56) /bd:[ Li0>D(20/56) Bi0>clk(16/61) Ro0<q(39/56) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input clk;    //: /sn:0 {0}(189,237)(215,237)(215,237)(257,237){1}
//: {2}(261,237)(311,237)(311,237)(378,237){3}
//: {4}(259,235)(259,172)(285,172){5}
output q;    //: /sn:0 {0}(558,185)(609,185)(609,185)(613,185){1}
input D;    //: /sn:0 {0}(291,93)(224,93)(224,149){1}
//: {2}(226,151)(272,151)(272,151)(285,151){3}
//: {4}(222,151)(185,151){5}
wire w7;    //: /sn:0 {0}(434,214)(444,214)(444,214)(491,214){1}
wire w4;    //: /sn:0 {0}(341,149)(462,149)(462,186)(491,186){1}
wire w10;    //: /sn:0 {0}(573,218)(558,218){1}
wire w2;    //: /sn:0 {0}(378,216)(359,216)(359,113)(333,113){1}
//: enddecls

  myAND g4 (.in0(clk), .in1(D), .out(w4));   //: @(286, 138) /sz:(54, 49) /R:1 /sn:0 /p:[ Li0>5 Li1>3 Ro0<0 ]
  //: joint g8 (clk) @(259, 237) /w:[ 2 4 1 -1 ]
  myINV g3 (.in(D), .out(w2));   //: @(292, 84) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  //: OUT g2 (q) @(610,185) /sn:0 /w:[ 1 ]
  //: IN g1 (clk) @(187,237) /sn:0 /w:[ 0 ]
  LatchSR g6 (.r(w7), .s(w4), .q(q), .nq(w10));   //: @(492, 164) /sz:(65, 76) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: joint g7 (D) @(224, 151) /w:[ 2 1 4 -1 ]
  myAND g5 (.in0(clk), .in1(w2), .out(w7));   //: @(379, 203) /sz:(54, 49) /R:1 /sn:0 /p:[ Li0>3 Li1>0 Ro0<0 ]
  //: IN g0 (D) @(183,151) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin myFA
module myFA(Cout, out, Cin, in1, in0);
//: interface  /sz:(54, 78) /bd:[ Ti0>in0(14/54) Ti1>in1(44/54) Li0>Cin(23/78) Bo0<out(25/54) Ro0<Cout(23/78) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(108,83)(137,83)(137,83)(139,83){1}
input Cin;    //: /sn:0 {0}(207,2)(207,26)(229,26){1}
input in0;    //: /sn:0 {0}(108,55)(139,55){1}
output out;    //: /sn:0 {0}(281,25)(326,25){1}
output Cout;    //: /sn:0 {0}(355,135)(386,135){1}
wire w0;    //: /sn:0 {0}(191,54)(229,54){1}
wire w8;    //: /sn:0 {0}(302,133)(175,133)(175,96){1}
wire w2;    //: /sn:0 {0}(265,67)(265,105)(302,105){1}
//: enddecls

  //: OUT g4 (Cout) @(383,135) /sn:0 /w:[ 1 ]
  //: OUT g3 (out) @(323,25) /sn:0 /w:[ 1 ]
  //: IN g2 (Cin) @(207,0) /sn:0 /R:3 /w:[ 0 ]
  //: IN g1 (in1) @(106,83) /sn:0 /w:[ 0 ]
  myHA g6 (.in1(w0), .in0(Cin), .Cout(w2), .out(out));   //: @(230, 17) /sz:(50, 49) /sn:0 /p:[ Li0>1 Li1>1 Bo0<0 Ro0<0 ]
  myOR g7 (.in0(w2), .in1(w8), .out(Cout));   //: @(303, 95) /sz:(51, 50) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  myHA g5 (.in1(in1), .in0(in0), .Cout(w8), .out(w0));   //: @(140, 46) /sz:(50, 49) /sn:0 /p:[ Li0>1 Li1>1 Bo0<1 Ro0<0 ]
  //: IN g0 (in0) @(106,55) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myCU
module myCU(c, enable, clk);
//: interface  /sz:(83, 55) /bd:[ Li0>enable(40/55) Li1>clk(14/55) Ro0<c(35/55) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input enable;    //: /sn:0 {0}(566,177)(566,222)(533,222){1}
input clk;    //: /sn:0 {0}(419,181)(419,247)(419,247)(419,290){1}
output c;    //: /sn:0 {0}(580,347)(580,345)(580,345)(580,380){1}
//: {2}(582,382)(619,382){3}
//: {4}(578,382)(445,382)(445,355){5}
wire w0;    //: /sn:0 {0}(449,290)(449,250)(474,250){1}
wire w1;    //: /sn:0 {0}(567,299)(567,251)(533,251){1}
//: enddecls

  myINV g4 (.in(c), .out(w1));   //: @(545, 300) /sz:(44, 46) /R:1 /sn:0 /p:[ Bi0>0 To0<0 ]
  FFDet g3 (.clk(clk), .D(w0), .q(c));   //: @(400, 291) /sz:(69, 63) /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<5 ]
  //: OUT g2 (c) @(616,382) /sn:0 /w:[ 3 ]
  //: IN g1 (enable) @(566,175) /sn:0 /R:3 /w:[ 0 ]
  //: joint g6 (c) @(580, 382) /w:[ 2 1 4 -1 ]
  myAND g5 (.in0(enable), .in1(w1), .out(w0));   //: @(475, 213) /sz:(57, 49) /R:3 /sn:0 /p:[ Ri0>1 Ri1>1 Lo0<1 ]
  //: IN g0 (clk) @(419,179) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNAND
module myNAND(out, in0, in1);
//: interface  /sz:(57, 58) /bd:[ Li0>in0(11/58) Li1>in1(44/58) Ro0<out(39/58) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w0;    //: /sn:0 {0}(100,49)(100,26)(134,26){1}
//: {2}(138,26)(171,26)(171,71){3}
//: {4}(136,24)(136,20)(136,20)(136,7){5}
input in1;    //: /sn:0 {0}(122,198)(47,198)(47,81){1}
//: {2}(49,79)(59,79)(59,79)(157,79){3}
//: {4}(45,79)(17,79){5}
supply0 w1;    //: /sn:0 {0}(136,207)(136,208)(136,208)(136,230){1}
input in0;    //: /sn:0 {0}(17,57)(67,57){1}
//: {2}(71,57)(84,57)(84,57)(86,57){3}
//: {4}(69,59)(69,145)(122,145){5}
output out;    //: /sn:0 {0}(136,137)(136,129)(136,129)(136,122){1}
//: {2}(138,120)(182,120)(182,120)(228,120){3}
//: {4}(136,118)(136,111)(136,111)(136,104){5}
//: {6}(138,102)(171,102)(171,88){7}
//: {8}(134,102)(100,102)(100,66){9}
wire w9;    //: /sn:0 {0}(136,154)(136,172)(136,172)(136,190){1}
//: enddecls

  //: OUT g8 (out) @(225,120) /sn:0 /w:[ 3 ]
  //: IN g4 (in0) @(15,57) /sn:0 /w:[ 0 ]
  //: joint g3 (out) @(136, 102) /w:[ 6 -1 8 5 ]
  _GGPMOS #(2, 1) pmos1 (.Z(out), .S(w0), .G(in1));   //: @(165,79) /w:[ 7 3 3 ]
  //: joint g2 (w0) @(136, 26) /w:[ 2 4 1 -1 ]
  //: GROUND g1 (w1) @(136,236) /sn:0 /w:[ 1 ]
  _GGNMOS #(2, 1) nmos1 (.Z(w9), .S(w1), .G(in1));   //: @(130,198) /w:[ 1 0 0 ]
  _GGNMOS #(2, 1) nmos0 (.Z(out), .S(w9), .G(in0));   //: @(130,145) /w:[ 0 0 5 ]
  //: joint g6 (in0) @(69, 57) /w:[ 2 -1 1 4 ]
  //: joint g9 (out) @(136, 120) /w:[ 2 4 -1 1 ]
  //: joint g7 (in1) @(47, 79) /w:[ 2 -1 4 1 ]
  //: IN g5 (in1) @(15,79) /sn:0 /w:[ 5 ]
  //: VDD g0 (w0) @(147,7) /sn:0 /w:[ 5 ]
  _GGPMOS #(2, 1) pmos0 (.Z(out), .S(w0), .G(in0));   //: @(94,57) /w:[ 9 0 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin LatchSR
module LatchSR(nq, q, r, s);
//: interface  /sz:(65, 76) /bd:[ Li0>r(50/76) Li1>s(22/76) Ro0<q(21/76) Ro1<nq(54/76) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input r;    //: /sn:0 {0}(78,203)(123,203){1}
output q;    //: /sn:0 {0}(123,176)(116,176)(116,136)(220,136)(220,113){1}
//: {2}(222,111)(262,111){3}
//: {4}(218,111)(178,111){5}
output nq;    //: /sn:0 {0}(181,203)(217,203){1}
//: {2}(221,203)(267,203){3}
//: {4}(219,201)(219,145)(98,145)(98,111)(120,111){5}
input s;    //: /sn:0 {0}(75,84)(107,84)(107,84)(120,84){1}
//: enddecls

  myNOR g4 (.in0(q), .in1(r), .out(nq));   //: @(124, 166) /sz:(56, 52) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 ]
  //: OUT g3 (nq) @(264,203) /sn:0 /w:[ 3 ]
  //: OUT g2 (q) @(259,111) /sn:0 /w:[ 3 ]
  //: IN g1 (r) @(76,203) /sn:0 /w:[ 0 ]
  //: joint g6 (q) @(220, 111) /w:[ 2 -1 4 1 ]
  //: joint g7 (nq) @(219, 203) /w:[ 2 4 1 -1 ]
  myNOR g5 (.in0(s), .in1(nq), .out(q));   //: @(121, 74) /sz:(56, 52) /sn:0 /p:[ Li0>1 Li1>5 Ro0<5 ]
  //: IN g0 (s) @(73,84) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin SQ4bit
module SQ4bit(out, in);
//: interface  /sz:(52, 59) /bd:[ Ti0>in[3:0](23/52) Bo0<out[7:0](26/52) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] in;    //: /sn:0 {0}(#:203,68)(233,68)(233,68)(238,68){1}
//: {2}(239,68)(276,68)(276,68)(293,68){3}
//: {4}(294,68)(335,68)(335,68)(376,68){5}
//: {6}(377,68)(415,68)(415,68)(452,68){7}
//: {8}(453,68)(482,68){9}
output [7:0] out;    //: /sn:0 {0}(#:632,708)(632,753){1}
supply0 w2;    //: /sn:0 {0}(586,666)(586,656)(607,656)(607,702){1}
wire w16;    //: /sn:0 {0}(570,182)(570,132)(503,132){1}
//: {2}(499,132)(404,132)(404,132)(322,132){3}
//: {4}(318,132)(300,132)(300,132)(296,132){5}
//: {6}(294,130)(294,92)(294,92)(294,72){7}
//: {8}(294,134)(294,149)(294,149)(294,181){9}
//: {10}(320,134)(320,228)(320,228)(320,322){11}
//: {12}(501,134)(501,144)(501,144)(501,182){13}
wire w6;    //: /sn:0 {0}(485,331)(485,286)(524,286)(524,238){1}
wire w7;    //: /sn:0 {0}(657,702)(657,634)(676,634)(676,563){1}
wire w4;    //: /sn:0 {0}(627,702)(627,626)(364,626)(364,447){1}
wire w3;    //: /sn:0 {0}(305,402)(305,640)(617,640)(617,702){1}
wire w0;    //: /sn:0 {0}(432,181)(432,155)(358,155){1}
//: {2}(354,155)(294,155)(294,155)(275,155){3}
//: {4}(271,155)(266,155)(266,155)(241,155){5}
//: {6}(239,153)(239,112)(239,112)(239,72){7}
//: {8}(239,157)(239,683)(597,683)(597,702){9}
//: {10}(273,157)(273,180)(273,180)(273,181){11}
//: {12}(356,157)(356,169)(356,169)(356,181){13}
wire w22;    //: /sn:0 {0}(706,507)(728,507)(728,663)(667,663)(667,702){1}
wire w20;    //: /sn:0 {0}(647,702)(647,601)(574,601)(574,563){1}
wire w30;    //: /sn:0 {0}(496,387)(563,387)(563,483){1}
wire w19;    //: /sn:0 {0}(496,356)(719,356)(719,115)(644,115){1}
//: {2}(640,115)(585,115)(585,115)(524,115){3}
//: {4}(520,115)(379,115){5}
//: {6}(377,113)(377,72){7}
//: {8}(377,117)(377,181){9}
//: {10}(522,117)(522,182){11}
//: {12}(642,117)(642,149)(642,149)(642,182){13}
wire w12;    //: /sn:0 {0}(298,322)(298,265)(298,265)(298,237){1}
wire w23;    //: /sn:0 {0}(593,238)(593,367)(593,367)(593,483){1}
wire w10;    //: /sn:0 {0}(637,702)(637,612)(451,612)(451,562){1}
wire w24;    //: /sn:0 {0}(665,483)(665,340)(665,340)(665,238){1}
wire w31;    //: /sn:0 {0}(432,508)(413,508)(413,392)(395,392){1}
wire w1;    //: /sn:0 {0}(359,367)(359,347)(336,347){1}
wire w32;    //: /sn:0 {0}(482,507)(491,507)(491,507)(548,507){1}
wire w8;    //: /sn:0 {0}(591,182)(591,100){1}
//: {2}(593,98)(630,98)(630,98)(661,98){3}
//: {4}(665,98)(733,98)(733,375)(695,375)(695,483){5}
//: {6}(663,100)(663,141)(663,141)(663,182){7}
//: {8}(589,98)(455,98){9}
//: {10}(453,96)(453,72){11}
//: {12}(453,100)(453,140)(453,140)(453,181){13}
wire w17;    //: /sn:0 {0}(604,507)(620,507)(620,507)(650,507){1}
wire w27;    //: /sn:0 {0}(466,482)(466,430)(466,430)(466,411){1}
wire w15;    //: /sn:0 {0}(379,367)(379,237){1}
wire w38;    //: /sn:0 {0}(455,331)(455,283)(455,283)(455,237){1}
//: enddecls

  myHA g8 (.in0(w12), .in1(w16), .out(w3), .Cout(w1));   //: @(287, 323) /sz:(48, 78) /sn:0 /p:[ Ti0>0 Ti1>11 Bo0<0 Ro0<1 ]
  //: joint g44 (w8) @(663, 98) /w:[ 4 -1 3 6 ]
  myAND g16 (.in1(w8), .in0(w0), .out(w38));   //: @(418, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>13 Ti1>0 Bo0<1 ]
  assign w0 = in[0]; //: TAP g3 @(239,66) /sn:0 /R:1 /w:[ 7 1 2 ] /ss:1
  //: joint g17 (w0) @(356, 155) /w:[ 1 -1 2 12 ]
  //: joint g26 (w8) @(453, 98) /w:[ 9 10 -1 12 ]
  assign out = {w22, w7, w20, w10, w4, w3, w2, w0}; //: CONCAT g2  @(632,707) /sn:0 /R:3 /w:[ 0 1 0 0 0 0 1 1 9 ] /dr:0 /tp:0 /drp:1
  //: comment g30 @(424,564) /sn:0
  //: /line:"HA3"
  //: /end
  //: joint g23 (w19) @(377, 115) /w:[ 5 6 -1 8 ]
  myAND g24 (.in1(w8), .in0(w19), .out(w24));   //: @(628, 183) /sz:(49, 54) /sn:0 /p:[ Ti0>7 Ti1>13 Bo0<1 ]
  //: OUT g1 (out) @(632,750) /sn:0 /R:3 /w:[ 1 ]
  //: comment g39 @(633,242) /sn:0
  //: /line:"a2a3"
  //: /end
  myHA g29 (.in1(w27), .in0(w31), .out(w10), .Cout(w32));   //: @(433, 483) /sz:(48, 78) /sn:0 /p:[ Ti0>0 Li0>0 Bo0<1 Ro0<0 ]
  myAND g18 (.in1(w19), .in0(w16), .out(w6));   //: @(487, 183) /sz:(49, 54) /sn:0 /p:[ Ti0>11 Ti1>13 Bo0<1 ]
  //: joint g10 (w0) @(239, 155) /w:[ 5 6 -1 8 ]
  //: joint g25 (w19) @(522, 115) /w:[ 3 -1 4 10 ]
  assign w19 = in[2]; //: TAP g6 @(377,66) /sn:0 /R:1 /w:[ 7 5 6 ] /ss:1
  myAND g9 (.in1(w16), .in0(w0), .out(w12));   //: @(259, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>9 Ti1>11 Bo0<1 ]
  assign w16 = in[1]; //: TAP g7 @(294,66) /sn:0 /R:1 /w:[ 7 3 4 ] /ss:1
  //: comment g35 @(439,414) /sn:0
  //: /line:"FA1"
  //: /end
  //: comment g31 @(260,383) /sn:0
  //: /line:"HA1"
  //: /end
  //: joint g22 (w16) @(501, 132) /w:[ 1 -1 2 12 ]
  //: comment g33 @(333,449) /sn:0
  //: /line:"HA2"
  //: /end
  //: comment g36 @(407,249) /sn:0
  //: /line:"a0a3"
  //: /end
  //: comment g41 @(546,566) /sn:0
  //: /line:"FA2"
  //: /end
  //: comment g42 @(650,565) /sn:0
  //: /line:"FA3"
  //: /end
  //: joint g40 (w19) @(642, 115) /w:[ 1 -1 2 12 ]
  myAND g12 (.in1(w19), .in0(w0), .out(w15));   //: @(342, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>9 Ti1>13 Bo0<1 ]
  myFA g28 (.in1(w6), .in0(w38), .Cin(w19), .out(w27), .Cout(w30));   //: @(441, 332) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Ro0<0 ]
  //: comment g34 @(340,241) /sn:0
  //: /line:"a0a2"
  //: /end
  myHA g14 (.in0(w1), .in1(w15), .out(w4), .Cout(w31));   //: @(346, 368) /sz:(48, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 Ro0<1 ]
  assign w8 = in[3]; //: TAP g5 @(453,66) /sn:0 /R:1 /w:[ 11 7 8 ] /ss:1
  //: joint g11 (w16) @(294, 132) /w:[ 5 6 -1 8 ]
  //: joint g19 (w16) @(320, 132) /w:[ 3 -1 4 10 ]
  myAND g21 (.in1(w8), .in0(w16), .out(w23));   //: @(556, 183) /sz:(49, 54) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  //: comment g32 @(259,242) /sn:0
  //: /line:"a0a1"
  //: /end
  //: GROUND ground (w2) @(586,672) /sn:0 /w:[ 0 ]
  myFA g15 (.in1(w8), .in0(w24), .Cin(w17), .out(w7), .Cout(w22));   //: @(651, 484) /sz:(54, 78) /sn:0 /p:[ Ti0>5 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  //: IN g0 (in) @(201,68) /sn:0 /w:[ 0 ]
  //: comment g38 @(559,239) /sn:0
  //: /line:"a1a3"
  //: /end
  //: joint g43 (w8) @(591, 98) /w:[ 2 -1 8 1 ]
  myFA g27 (.in1(w23), .in0(w30), .Cin(w32), .out(w20), .Cout(w17));   //: @(549, 484) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  //: comment g37 @(491,243) /sn:0
  //: /line:"a1a2"
  //: /end
  //: joint g13 (w0) @(273, 155) /w:[ 3 -1 4 10 ]

endmodule
//: /netlistEnd

//: /netlistBegin myEXOR
module myEXOR(out, in1, in0);
//: interface  /sz:(52, 55) /bd:[ Li0>in1(44/55) Li1>in0(12/55) Ro0<out(42/55) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(198,81)(80,81)(80,140){1}
//: {2}(82,142)(94,142){3}
//: {4}(78,142)(69,142)(69,142)(57,142){5}
input in0;    //: /sn:0 {0}(198,129)(166,129)(166,70)(82,70){1}
//: {2}(80,68)(80,28)(95,28){3}
//: {4}(78,70)(54,70){5}
output out;    //: /sn:0 {0}(357,130)(384,130)(384,130)(387,130){1}
wire w6;    //: /sn:0 {0}(257,76)(278,76)(278,102)(298,102){1}
wire w3;    //: /sn:0 {0}(136,162)(107,162)(107,162)(198,162){1}
wire w1;    //: /sn:0 {0}(137,48)(107,48)(107,48)(198,48){1}
wire w9;    //: /sn:0 {0}(257,157)(278,157)(278,135)(298,135){1}
//: enddecls

  myINV g4 (.in(in1), .out(w3));   //: @(95, 133) /sz:(40, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  myNAND g8 (.in0(in0), .in1(w3), .out(w9));   //: @(199, 118) /sz:(57, 58) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 ]
  myINV g3 (.in(in0), .out(w1));   //: @(96, 19) /sz:(40, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: OUT g2 (out) @(384,130) /sn:0 /w:[ 1 ]
  //: IN g1 (in1) @(55,142) /sn:0 /w:[ 5 ]
  //: joint g6 (in0) @(80, 70) /w:[ 1 2 4 -1 ]
  myNAND g7 (.in0(w6), .in1(w9), .out(out));   //: @(299, 91) /sz:(57, 58) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: joint g9 (in1) @(80, 142) /w:[ 2 1 4 -1 ]
  myNAND g5 (.in0(w1), .in1(in1), .out(w6));   //: @(199, 37) /sz:(57, 58) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  //: IN g0 (in0) @(52,70) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUL4x4
module MUL4x4(b, p, a);
//: interface  /sz:(65, 59) /bd:[ Ti0>a[3:0](18/65) Ti1>b[3:0](41/65) Bo0<p[7:0](32/65) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output [7:0] p;    //: /sn:0 {0}(527,817)(#:527,774){1}
input [3:0] b;    //: /sn:0 {0}(#:883,136)(875,136){1}
//: {2}(874,136)(648,136){3}
//: {4}(647,136)(419,136){5}
//: {6}(418,136)(193,136){7}
//: {8}(192,136)(#:133,136){9}
input [3:0] a;    //: /sn:0 {0}(#:133,48)(171,48){1}
//: {2}(172,48)(227,48){3}
//: {4}(228,48)(283,48){5}
//: {6}(284,48)(340,48){7}
//: {8}(341,48)(347,48){9}
wire w16;    //: /sn:0 {0}(532,768)(532,719)(598,719)(598,694){1}
wire w13;    //: /sn:0 {0}(512,768)(512,727)(360,727)(360,553){1}
wire w6;    //: /sn:0 {0}(970,181)(970,86)(742,86){1}
//: {2}(738,86)(513,86){3}
//: {4}(509,86)(286,86){5}
//: {6}(284,84)(284,62)(284,62)(284,52){7}
//: {8}(284,88)(284,181){9}
//: {10}(511,88)(511,134)(511,134)(511,181){11}
//: {12}(740,88)(740,181){13}
wire w7;    //: /sn:0 {0}(258,405)(258,737)(502,737)(502,768){1}
wire w50;    //: /sn:0 {0}(862,350)(919,350)(919,615){1}
wire w34;    //: /sn:0 {0}(484,350)(545,350)(545,350)(567,350){1}
wire w39;    //: /sn:0 {0}(623,350)(723,350)(723,350)(806,350){1}
wire w4;    //: /sn:0 {0}(912,181)(912,101)(685,101){1}
//: {2}(681,101)(457,101){3}
//: {4}(453,101)(230,101){5}
//: {6}(228,99)(228,70)(228,70)(228,52){7}
//: {8}(228,103)(228,181){9}
//: {10}(455,103)(455,181){11}
//: {12}(683,103)(683,181){13}
wire w36;    //: /sn:0 {0}(593,474)(593,429)(593,429)(593,406){1}
wire w22;    //: /sn:0 {0}(289,350)(327,350){1}
wire w0;    //: /sn:0 {0}(362,181)(362,163)(307,163){1}
//: {2}(303,163)(251,163){3}
//: {4}(247,163)(195,163){5}
//: {6}(193,161)(193,140){7}
//: {8}(193,165)(193,181){9}
//: {10}(249,165)(249,181){11}
//: {12}(305,165)(305,181){13}
wire w20;    //: /sn:0 {0}(534,237)(534,291)(473,291)(473,326){1}
wire w30;    //: /sn:0 {0}(1049,237)(1049,370)(949,370)(949,615){1}
wire w29;    //: /sn:0 {0}(706,237)(706,448)(484,448)(484,474){1}
wire w42;    //: /sn:0 {0}(465,614)(465,593)(465,593)(465,554){1}
wire w37;    //: /sn:0 {0}(1047,181)(1047,164)(993,164){1}
//: {2}(989,164)(935,164){3}
//: {4}(931,164)(877,164){5}
//: {6}(875,162)(875,140){7}
//: {8}(875,166)(875,181){9}
//: {10}(933,166)(933,181){11}
//: {12}(991,166)(991,181){13}
wire w19;    //: /sn:0 {0}(918,695)(918,740)(552,740)(552,768){1}
wire w18;    //: /sn:0 {0}(813,695)(813,728)(542,728)(542,768){1}
wire w12;    //: /sn:0 {0}(590,181)(590,164)(534,164){1}
//: {2}(530,164)(478,164){3}
//: {4}(474,164)(421,164){5}
//: {6}(419,162)(419,140){7}
//: {8}(419,166)(419,181){9}
//: {10}(476,166)(476,181){11}
//: {12}(532,166)(532,173)(532,173)(532,181){13}
wire w23;    //: /sn:0 {0}(592,237)(592,264)(582,264)(582,326){1}
wire w21;    //: /sn:0 {0}(562,768)(562,758)(970,758)(970,669)(960,669){1}
wire w24;    //: /sn:0 {0}(819,181)(819,162)(763,162){1}
//: {2}(759,162)(706,162){3}
//: {4}(702,162)(650,162){5}
//: {6}(648,160)(648,140){7}
//: {8}(648,164)(648,181){9}
//: {10}(704,164)(704,181){11}
//: {12}(761,164)(761,181){13}
wire w31;    //: /sn:0 {0}(503,639)(575,639){1}
wire w1;    //: /sn:0 {0}(854,181)(854,120)(629,120){1}
//: {2}(625,120)(400,120){3}
//: {4}(396,120)(174,120){5}
//: {6}(172,118)(172,79)(172,79)(172,52){7}
//: {8}(172,122)(172,181){9}
//: {10}(398,122)(398,181){11}
//: {12}(627,122)(627,181){13}
wire w32;    //: /sn:0 {0}(821,237)(821,297)(821,297)(821,326){1}
wire w46;    //: /sn:0 {0}(634,498)(802,498)(802,615){1}
wire w8;    //: /sn:0 {0}(307,237)(307,311)(342,311)(342,326){1}
wire w52;    //: /sn:0 {0}(843,639)(882,639)(882,639)(904,639){1}
wire w27;    //: /sn:0 {0}(353,473)(353,406){1}
wire w17;    //: /sn:0 {0}(478,237)(478,280)(372,280)(372,326){1}
wire w44;    //: /sn:0 {0}(935,237)(935,459)(623,459)(623,474){1}
wire w33;    //: /sn:0 {0}(454,406)(454,474){1}
wire w28;    //: /sn:0 {0}(383,350)(428,350){1}
wire w35;    //: /sn:0 {0}(763,237)(763,281)(612,281)(612,326){1}
wire w49;    //: /sn:0 {0}(832,406)(832,510)(832,510)(832,615){1}
wire w45;    //: /sn:0 {0}(604,614)(604,588)(604,588)(604,554){1}
wire w14;    //: /sn:0 {0}(273,325)(273,273)(421,273)(421,237){1}
wire w48;    //: /sn:0 {0}(634,639)(719,639)(719,639)(787,639){1}
wire w2;    //: /sn:0 {0}(492,768)(492,747)(195,747)(195,237){1}
wire w11;    //: /sn:0 {0}(364,237)(364,301)(443,301)(443,326){1}
wire w41;    //: /sn:0 {0}(993,237)(993,311)(851,311)(851,326){1}
wire w15;    //: /sn:0 {0}(472,694)(472,719)(522,719)(522,768){1}
wire w5;    //: /sn:0 {0}(251,325)(251,237){1}
wire w38;    //: /sn:0 {0}(877,237)(877,595)(487,595)(487,614){1}
wire w43;    //: /sn:0 {0}(495,498)(556,498)(556,498)(578,498){1}
wire w9;    //: /sn:0 {0}(1026,181)(1026,70)(800,70){1}
//: {2}(796,70)(571,70){3}
//: {4}(567,70)(343,70){5}
//: {6}(341,68)(341,52){7}
//: {8}(341,72)(341,181){9}
//: {10}(569,72)(569,181){11}
//: {12}(798,72)(798,181){13}
wire w26;    //: /sn:0 {0}(650,237)(650,436)(375,436)(375,473){1}
wire w40;    //: /sn:0 {0}(391,498)(418,498)(418,498)(439,498){1}
//: enddecls

  myAND g4 (.in0(w1), .in1(w12), .out(w14));   //: @(384, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>11 Ti1>9 Bo0<1 ]
  myAND g8 (.in0(w6), .in1(w12), .out(w20));   //: @(497, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>11 Ti1>13 Bo0<0 ]
  //: joint g44 (w4) @(683, 101) /w:[ 1 -1 2 12 ]
  myAND g3 (.in0(w4), .in1(w0), .out(w5));   //: @(214, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>9 Ti1>11 Bo0<1 ]
  myAND g16 (.in0(w6), .in1(w37), .out(w41));   //: @(956, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>0 Ti1>13 Bo0<0 ]
  //: joint g47 (w37) @(875, 164) /w:[ 5 6 -1 8 ]
  myAND g17 (.in0(w4), .in1(w37), .out(w44));   //: @(898, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>0 Ti1>11 Bo0<0 ]
  assign w12 = b[1]; //: TAP g26 @(419,134) /sn:0 /R:1 /w:[ 7 6 5 ] /ss:1
  myAND g2 (.in0(w1), .in1(w0), .out(w2));   //: @(158, 182) /sz:(49, 54) /R:3 /sn:0 /p:[ Ti0>9 Ti1>9 Bo0<1 ]
  //: joint g23 (w0) @(249, 163) /w:[ 3 -1 4 10 ]
  //: joint g30 (w9) @(341, 70) /w:[ 5 6 -1 8 ]
  //: IN g1 (b) @(131,136) /sn:0 /w:[ 9 ]
  //: joint g24 (w0) @(305, 163) /w:[ 1 -1 2 12 ]
  //: joint g39 (w4) @(455, 101) /w:[ 3 -1 4 10 ]
  myHA g60 (.in1(w45), .in0(w31), .out(w16), .Cout(w48));   //: @(576, 615) /sz:(57, 78) /sn:0 /p:[ Ti0>0 Li0>1 Bo0<1 Ro0<0 ]
  //: joint g29 (w6) @(284, 86) /w:[ 5 6 -1 8 ]
  assign p = {w21, w19, w18, w16, w15, w13, w7, w2}; //: CONCAT g51  @(527,773) /sn:0 /R:3 /w:[ 1 0 1 1 0 1 0 1 0 ] /dr:0 /tp:0 /drp:1
  myAND g18 (.in0(w9), .in1(w37), .out(w30));   //: @(1012, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  myAND g10 (.in0(w1), .in1(w24), .out(w26));   //: @(613, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>13 Ti1>9 Bo0<0 ]
  assign w9 = a[3]; //: TAP g25 @(341,46) /sn:0 /R:1 /w:[ 7 7 8 ] /ss:1
  //: joint g49 (w37) @(991, 164) /w:[ 1 -1 2 12 ]
  myAND g6 (.in0(w9), .in1(w0), .out(w11));   //: @(327, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>9 Ti1>0 Bo0<0 ]
  //: OUT g50 (p) @(527,814) /sn:0 /R:3 /w:[ 0 ]
  myFA g58 (.in1(w35), .in0(w23), .Cin(w34), .out(w36), .Cout(w39));   //: @(568, 327) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  myFA g56 (.in1(w29), .in0(w33), .Cin(w40), .out(w42), .Cout(w43));   //: @(440, 475) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  myAND g7 (.in0(w4), .in1(w12), .out(w17));   //: @(441, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>11 Ti1>11 Bo0<0 ]
  myAND g9 (.in0(w9), .in1(w12), .out(w23));   //: @(555, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>11 Ti1>0 Bo0<0 ]
  assign w24 = b[2]; //: TAP g35 @(648,134) /sn:0 /R:1 /w:[ 7 4 3 ] /ss:1
  myFA g59 (.in1(w44), .in0(w36), .Cin(w43), .out(w45), .Cout(w46));   //: @(579, 475) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  assign w6 = a[2]; //: TAP g22 @(284,46) /sn:0 /R:1 /w:[ 7 5 6 ] /ss:1
  //: joint g31 (w12) @(419, 164) /w:[ 5 6 -1 8 ]
  myFA g54 (.in1(w20), .in0(w11), .Cin(w28), .out(w33), .Cout(w34));   //: @(429, 327) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  //: joint g33 (w12) @(532, 164) /w:[ 1 -1 2 12 ]
  //: joint g36 (w24) @(648, 162) /w:[ 5 6 -1 8 ]
  //: joint g41 (w9) @(569, 70) /w:[ 3 -1 4 10 ]
  //: joint g45 (w6) @(740, 86) /w:[ 1 -1 2 12 ]
  myHA g52 (.in0(w5), .in1(w14), .out(w7), .Cout(w22));   //: @(240, 326) /sz:(48, 78) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Ro0<0 ]
  //: joint g40 (w6) @(511, 86) /w:[ 3 -1 4 10 ]
  //: joint g42 (w1) @(627, 120) /w:[ 1 -1 2 12 ]
  assign w1 = a[0]; //: TAP g12 @(172,46) /sn:0 /R:1 /w:[ 7 1 2 ] /ss:1
  myHA g57 (.in0(w42), .in1(w38), .out(w15), .Cout(w31));   //: @(454, 615) /sz:(48, 78) /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<0 Ro0<0 ]
  //: joint g28 (w4) @(228, 101) /w:[ 5 6 -1 8 ]
  //: joint g34 (w1) @(398, 120) /w:[ 3 -1 4 10 ]
  //: joint g46 (w9) @(798, 70) /w:[ 1 -1 2 12 ]
  myAND g5 (.in0(w6), .in1(w0), .out(w8));   //: @(270, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>9 Ti1>13 Bo0<0 ]
  myAND g11 (.in0(w4), .in1(w24), .out(w29));   //: @(669, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>13 Ti1>11 Bo0<0 ]
  myAND g14 (.in0(w6), .in1(w24), .out(w35));   //: @(726, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>13 Ti1>13 Bo0<0 ]
  myFA g61 (.in1(w41), .in0(w32), .Cin(w39), .out(w49), .Cout(w50));   //: @(807, 327) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  assign w0 = b[0]; //: TAP g19 @(193,134) /sn:0 /R:1 /w:[ 7 8 7 ] /ss:1
  //: joint g21 (w0) @(193, 163) /w:[ 5 6 -1 8 ]
  assign w4 = a[1]; //: TAP g20 @(228,46) /sn:0 /R:1 /w:[ 7 3 4 ] /ss:1
  //: joint g32 (w12) @(476, 164) /w:[ 3 -1 4 10 ]
  myFA g63 (.in1(w30), .in0(w50), .Cin(w52), .out(w19), .Cout(w21));   //: @(905, 616) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<1 ]
  //: IN g0 (a) @(131,48) /sn:0 /w:[ 0 ]
  myAND g15 (.in0(w1), .in1(w37), .out(w38));   //: @(840, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>0 Ti1>9 Bo0<0 ]
  //: joint g38 (w24) @(761, 162) /w:[ 1 -1 2 12 ]
  assign w37 = b[3]; //: TAP g43 @(875,134) /sn:0 /R:1 /w:[ 7 2 1 ] /ss:1
  //: joint g27 (w1) @(172, 120) /w:[ 5 6 -1 8 ]
  //: joint g48 (w37) @(933, 164) /w:[ 3 -1 4 10 ]
  myFA g62 (.in1(w49), .in0(w46), .Cin(w48), .out(w18), .Cout(w52));   //: @(788, 616) /sz:(54, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  //: joint g37 (w24) @(704, 162) /w:[ 3 -1 4 10 ]
  myHA g55 (.in0(w27), .in1(w26), .out(w13), .Cout(w40));   //: @(342, 474) /sz:(48, 78) /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<1 Ro0<0 ]
  myFA g53 (.in1(w17), .in0(w8), .Cin(w22), .out(w27), .Cout(w28));   //: @(328, 327) /sz:(54, 78) /R:2 /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]
  myAND g13 (.in0(w9), .in1(w24), .out(w32));   //: @(784, 182) /sz:(49, 54) /sn:0 /p:[ Ti0>13 Ti1>0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDet
module FFDet(q, clk, D);
//: interface  /sz:(69, 63) /bd:[ Ti0>clk(54/69) Ti1>D(17/69) Bo0<q(45/69) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input clk;    //: /sn:0 {0}(250,267)(213,267){1}
//: {2}(209,267)(182,267){3}
//: {4}(211,269)(211,343)(429,343)(429,333){5}
output q;    //: /sn:0 {0}(475,315)(529,315){1}
input D;    //: /sn:0 {0}(183,200)(246,200)(246,200)(305,200){1}
wire w1;    //: /sn:0 {0}(292,287)(322,287)(322,237){1}
wire w2;    //: /sn:0 {0}(368,219)(392,219)(392,296)(412,296){1}
//: enddecls

  FFDls g4 (.D(w2), .clk(clk), .q(q));   //: @(413, 276) /sz:(61, 56) /sn:0 /p:[ Li0>1 Bi0>5 Ro0<0 ]
  FFDls g3 (.D(D), .clk(w1), .q(w2));   //: @(306, 180) /sz:(61, 56) /sn:0 /p:[ Li0>1 Bi0>1 Ro0<0 ]
  //: OUT g2 (q) @(526,315) /sn:0 /w:[ 1 ]
  //: IN g1 (clk) @(180,267) /sn:0 /w:[ 3 ]
  //: joint g6 (clk) @(211, 267) /w:[ 1 -1 2 4 ]
  myINV g5 (.in(clk), .out(w1));   //: @(251, 258) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: IN g0 (D) @(181,200) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX4bit
module MUX4bit(out, c, b, a);
//: interface  /sz:(68, 64) /bd:[ Ti0>b[3:0](44/68) Ti1>a[3:0](17/68) Li0>c(35/64) Bo0<out[3:0](31/68) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:299,92)(400,92){1}
//: {2}(401,92)(445,92)(445,92)(488,92){3}
//: {4}(489,92)(577,92){5}
//: {6}(578,92)(668,92){7}
//: {8}(669,92)(680,92){9}
output [3:0] out;    //: /sn:0 {0}(526,304)(#:526,271){1}
input [3:0] a;    //: /sn:0 {0}(#:297,59)(374,59){1}
//: {2}(375,59)(419,59)(419,59)(462,59){3}
//: {4}(463,59)(551,59){5}
//: {6}(552,59)(597,59)(597,59)(642,59){7}
//: {8}(643,59)(652,59){9}
input c;    //: /sn:0 {0}(298,131)(319,131)(319,131)(343,131){1}
//: {2}(347,131)(386,131)(386,131)(434,131){3}
//: {4}(438,131)(468,131)(468,131)(521,131){5}
//: {6}(525,131)(617,131)(617,176)(627,176){7}
//: {8}(523,133)(523,177)(536,177){9}
//: {10}(436,133)(436,177)(447,177){11}
//: {12}(345,133)(345,178)(359,178){13}
wire w13;    //: /sn:0 {0}(401,96)(401,137)(401,137)(401,156){1}
wire w7;    //: /sn:0 {0}(541,265)(541,243)(656,243)(656,201){1}
wire w4;    //: /sn:0 {0}(643,63)(643,123)(643,123)(643,154){1}
wire w3;    //: /sn:0 {0}(531,265)(531,233)(567,233)(567,202){1}
wire w0;    //: /sn:0 {0}(552,63)(552,124)(552,124)(552,155){1}
wire w12;    //: /sn:0 {0}(375,63)(375,124)(375,124)(375,156){1}
wire w1;    //: /sn:0 {0}(578,96)(578,136)(578,136)(578,155){1}
wire w8;    //: /sn:0 {0}(463,63)(463,124)(463,124)(463,155){1}
wire w11;    //: /sn:0 {0}(521,265)(521,232)(477,232)(477,202){1}
wire w15;    //: /sn:0 {0}(389,203)(389,244)(511,244)(511,265){1}
wire w5;    //: /sn:0 {0}(669,96)(669,136)(669,136)(669,154){1}
wire w9;    //: /sn:0 {0}(489,96)(489,136)(489,136)(489,155){1}
//: enddecls

  //: joint g8 (c) @(523, 131) /w:[ 6 -1 5 8 ]
  MUX g4 (.b(w1), .a(w0), .c(c), .out(w3));   //: @(537, 156) /sz:(56, 45) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>9 Bo0<1 ]
  assign w8 = a[1]; //: TAP g16 @(463,57) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: OUT g3 (out) @(526,301) /sn:0 /R:3 /w:[ 0 ]
  assign w13 = b[0]; //: TAP g17 @(401,90) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: IN g2 (c) @(296,131) /sn:0 /w:[ 0 ]
  //: IN g1 (b) @(297,92) /sn:0 /w:[ 0 ]
  assign w12 = a[0]; //: TAP g18 @(375,57) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g10 (c) @(345, 131) /w:[ 2 -1 1 12 ]
  MUX g6 (.b(w9), .a(w8), .c(c), .out(w11));   //: @(448, 156) /sz:(56, 45) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>11 Bo0<1 ]
  //: joint g9 (c) @(436, 131) /w:[ 4 -1 3 10 ]
  MUX g7 (.b(w13), .a(w12), .c(c), .out(w15));   //: @(360, 157) /sz:(56, 45) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>13 Bo0<0 ]
  assign w4 = a[3]; //: TAP g12 @(643,57) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w0 = a[2]; //: TAP g14 @(552,57) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w5 = b[3]; //: TAP g11 @(669,90) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  MUX g5 (.b(w5), .a(w4), .c(c), .out(w7));   //: @(628, 155) /sz:(56, 45) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Li0>7 Bo0<1 ]
  assign out = {w7, w3, w11, w15}; //: CONCAT g19  @(526,270) /sn:0 /R:3 /w:[ 1 0 0 0 1 ] /dr:0 /tp:0 /drp:1
  assign w9 = b[1]; //: TAP g15 @(489,90) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: IN g0 (a) @(295,59) /sn:0 /w:[ 0 ]
  assign w1 = b[2]; //: TAP g13 @(578,90) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin myOR
module myOR(out, in1, in0);
//: interface  /sz:(51, 50) /bd:[ Li0>in0(10/50) Li1>in1(38/50) Ro0<out(40/50) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(64,96)(86,96)(86,96)(102,96){1}
input in0;    //: /sn:0 {0}(64,69)(87,69)(87,69)(102,69){1}
output out;    //: /sn:0 {0}(235,116)(245,116)(245,116)(269,116){1}
wire w2;    //: /sn:0 {0}(160,96)(178,96)(178,96)(193,96){1}
//: enddecls

  //: OUT g4 (out) @(266,116) /sn:0 /w:[ 1 ]
  myINV g3 (.in(w2), .out(out));   //: @(194, 87) /sz:(40, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  myNOR g2 (.in1(in1), .in0(in0), .out(w2));   //: @(103, 59) /sz:(56, 52) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g1 (in1) @(62,96) /sn:0 /w:[ 0 ]
  //: IN g0 (in0) @(62,69) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNOR
module myNOR(out, in1, in0);
//: interface  /sz:(56, 52) /bd:[ Li0>in0(10/52) Li1>in1(37/52) Ro0<out(37/52) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w0;    //: /sn:0 {0}(161,12)(161,29)(161,29)(161,41){1}
input in1;    //: /sn:0 {0}(52,107)(116,107)(116,107)(130,107){1}
//: {2}(134,107)(147,107){3}
//: {4}(132,109)(132,199)(179,199){5}
supply0 w1;    //: /sn:0 {0}(115,235)(115,248)(163,248){1}
//: {2}(167,248)(193,248)(193,208){3}
//: {4}(165,250)(165,244)(165,244)(165,268){5}
input in0;    //: /sn:0 {0}(50,49)(65,49)(65,49)(80,49){1}
//: {2}(84,49)(115,49)(115,49)(147,49){3}
//: {4}(82,51)(82,226)(101,226){5}
output out;    //: /sn:0 {0}(193,191)(193,173)(163,173){1}
//: {2}(161,171)(161,145){3}
//: {4}(163,143)(93,143)(93,143)(233,143){5}
//: {6}(161,141)(161,116){7}
//: {8}(159,173)(115,173)(115,218){9}
wire w2;    //: /sn:0 {0}(161,58)(161,78)(161,78)(161,99){1}
//: enddecls

  //: joint g8 (in0) @(82, 49) /w:[ 2 -1 1 4 ]
  //: GROUND g4 (w1) @(165,274) /sn:0 /w:[ 5 ]
  _GGPMOS #(2, 1) pmos1 (.Z(out), .S(w2), .G(in1));   //: @(155,107) /w:[ 7 1 3 ]
  //: VDD g3 (w0) @(172,12) /sn:0 /w:[ 0 ]
  //: OUT g2 (out) @(230,143) /sn:0 /w:[ 5 ]
  //: IN g1 (in1) @(50,107) /sn:0 /w:[ 0 ]
  _GGNMOS #(2, 1) nmos1 (.Z(out), .S(w1), .G(in1));   //: @(187,199) /w:[ 0 3 5 ]
  _GGNMOS #(2, 1) nmos0 (.Z(out), .S(w1), .G(in0));   //: @(109,226) /w:[ 9 0 5 ]
  //: joint g6 (out) @(161, 143) /w:[ 4 6 -1 3 ]
  //: joint g9 (in1) @(132, 107) /w:[ 2 -1 1 4 ]
  //: joint g7 (w1) @(165, 248) /w:[ 2 -1 1 4 ]
  //: joint g5 (out) @(161, 173) /w:[ 1 2 8 -1 ]
  //: IN g0 (in0) @(48,49) /sn:0 /w:[ 0 ]
  _GGPMOS #(2, 1) pmos0 (.Z(w2), .S(w0), .G(in0));   //: @(155,49) /w:[ 0 1 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin myAND
module myAND(out, in1, in0);
//: interface  /sz:(49, 54) /bd:[ Ti0>in0(14/49) Ti1>in1(35/49) Bo0<out(37/49) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(101,135)(131,135)(131,135)(146,135){1}
input in0;    //: /sn:0 {0}(103,102)(131,102)(131,102)(146,102){1}
output out;    //: /sn:0 {0}(290,150)(321,150)(321,150)(324,150){1}
wire w2;    //: /sn:0 {0}(205,130)(233,130)(233,130)(248,130){1}
//: enddecls

  //: OUT g4 (out) @(321,150) /sn:0 /w:[ 1 ]
  myINV g3 (.in(w2), .out(out));   //: @(249, 121) /sz:(40, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  myNAND g2 (.in1(in1), .in0(in0), .out(w2));   //: @(147, 91) /sz:(57, 58) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g1 (in1) @(99,135) /sn:0 /w:[ 0 ]
  //: IN g0 (in0) @(101,102) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myINV
module myINV(in, out);
//: interface  /sz:(40, 40) /bd:[ Li0>in(9/40) Ro0<out(29/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in;    //: /sn:0 {0}(181,133)(146,133)(146,96){1}
//: {2}(148,94)(154,94)(154,94)(122,94){3}
//: {4}(146,92)(146,59)(181,59){5}
supply1 w0;    //: /sn:0 {0}(195,51)(195,11){1}
supply0 w1;    //: /sn:0 {0}(195,173)(195,142){1}
output out;    //: /sn:0 {0}(195,125)(195,96){1}
//: {2}(197,94)(226,94)(226,94)(230,94){3}
//: {4}(195,92)(195,68){5}
//: enddecls

  //: IN g4 (in) @(120,94) /sn:0 /w:[ 3 ]
  //: GROUND g1 (w1) @(195,179) /sn:0 /w:[ 0 ]
  _GGNMOS #(2, 1) nmos0 (.Z(out), .S(w1), .G(in));   //: @(189,133) /w:[ 0 1 0 ]
  //: OUT g6 (out) @(227,94) /sn:0 /w:[ 3 ]
  //: joint g7 (out) @(195, 94) /w:[ 2 4 -1 1 ]
  //: joint g5 (in) @(146, 94) /w:[ 2 4 -1 1 ]
  //: VDD g0 (w0) @(206,11) /sn:0 /w:[ 1 ]
  _GGPMOS #(2, 1) pmos0 (.Z(out), .S(w0), .G(in));   //: @(189,59) /w:[ 5 0 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX
module MUX(out, c, b, a);
//: interface  /sz:(56, 45) /bd:[ Ti0>a(15/56) Ti1>b(41/56) Li0>c(21/45) Bo0<out(36/56) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(246,315)(304,315)(304,315)(379,315){1}
output out;    //: /sn:0 {0}(550,271)(597,271){1}
input a;    //: /sn:0 {0}(244,184)(307,184)(307,184)(380,184){1}
input c;    //: /sn:0 {0}(379,282)(266,282)(266,240){1}
//: {2}(268,238)(299,238){3}
//: {4}(264,238)(263,238)(263,238)(245,238){5}
wire w7;    //: /sn:0 {0}(438,310)(468,310)(468,276)(491,276){1}
wire w4;    //: /sn:0 {0}(439,212)(467,212)(467,243)(491,243){1}
wire w1;    //: /sn:0 {0}(341,217)(373,217)(373,217)(380,217){1}
//: enddecls

  //: joint g8 (c) @(266, 238) /w:[ 2 -1 4 1 ]
  myINV g4 (.in(c), .out(w1));   //: @(300, 209) /sz:(40, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: OUT g3 (out) @(594,271) /sn:0 /w:[ 1 ]
  //: IN g2 (c) @(243,238) /sn:0 /w:[ 5 ]
  //: IN g1 (b) @(244,315) /sn:0 /w:[ 0 ]
  myNAND g6 (.in1(b), .in0(c), .out(w7));   //: @(380, 271) /sz:(57, 58) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  myNAND g7 (.in1(w7), .in0(w4), .out(out));   //: @(492, 232) /sz:(57, 58) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  myNAND g5 (.in1(w1), .in0(a), .out(w4));   //: @(381, 173) /sz:(57, 58) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g0 (a) @(242,184) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin RCA8bit
module RCA8bit(out, b, C0, a);
//: interface  /sz:(67, 75) /bd:[ Li0>b[7:0](61/75) Li1>a[7:0](12/75) Ro0<out[8:0](47/75) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] b;    //: /sn:0 {0}(#:978,196)(963,196){1}
//: {2}(962,196)(920,196)(920,196)(877,196){3}
//: {4}(876,196)(786,196){5}
//: {6}(785,196)(742,196)(742,196)(698,196){7}
//: {8}(697,196)(611,196){9}
//: {10}(610,196)(523,196){11}
//: {12}(522,196)(435,196){13}
//: {14}(434,196)(348,196){15}
//: {16}(347,196)(#:253,196){17}
input C0;    //: {0}(303,256)(280,256)(280,256)(99:254,256){1}
output [8:0] out;    //: /sn:0 {0}(679,487)(679,434)(#:679,434)(#:679,439){1}
input [7:0] a;    //: /sn:0 {0}(#:985,166)(933,166){1}
//: {2}(932,166)(890,166)(890,166)(847,166){3}
//: {4}(846,166)(756,166){5}
//: {6}(755,166)(668,166){7}
//: {8}(667,166)(581,166){9}
//: {10}(580,166)(493,166){11}
//: {12}(492,166)(405,166){13}
//: {14}(404,166)(318,166){15}
//: {16}(317,166)(#:252,166){17}
wire w13;    //: /sn:0 {0}(709,433)(709,392)(944,392)(944,312){1}
wire w6;    //: /sn:0 {0}(649,433)(649,390)(416,390)(416,312){1}
wire w16;    //: /sn:0 {0}(405,232)(405,170){1}
wire w34;    //: /sn:0 {0}(756,232)(756,170){1}
wire w39;    //: /sn:0 {0}(847,232)(847,178)(847,178)(847,170){1}
wire w25;    //: /sn:0 {0}(611,232)(611,200){1}
wire w4;    //: /sn:0 {0}(359,256)(375,256)(375,256)(390,256){1}
wire w3;    //: /sn:0 {0}(639,433)(639,406)(329,406)(329,312){1}
wire w0;    //: /sn:0 {0}(318,232)(318,170){1}
wire w20;    //: /sn:0 {0}(523,232)(523,200){1}
wire w30;    //: /sn:0 {0}(698,232)(698,208)(698,208)(698,200){1}
wire w19;    //: /sn:0 {0}(493,232)(493,170){1}
wire w18;    //: /sn:0 {0}(446,256)(460,256)(460,256)(478,256){1}
wire w12;    //: /sn:0 {0}(699,433)(699,380)(858,380)(858,312){1}
wire w23;    //: /sn:0 {0}(534,256)(533,256)(533,256)(566,256){1}
wire w10;    //: /sn:0 {0}(679,433)(679,372)(679,372)(679,312){1}
wire w1;    //: /sn:0 {0}(348,232)(348,200){1}
wire w8;    //: /sn:0 {0}(659,433)(659,380)(504,380)(504,312){1}
wire w44;    //: /sn:0 {0}(933,232)(933,178)(933,178)(933,170){1}
wire w17;    //: /sn:0 {0}(668,232)(668,170){1}
wire w35;    //: /sn:0 {0}(786,232)(786,200){1}
wire w33;    //: /sn:0 {0}(741,256)(716,256)(716,258)(716,258)(716,256)(709,256){1}
wire w28;    //: /sn:0 {0}(622,256)(624,256)(624,256)(653,256){1}
wire w45;    //: /sn:0 {0}(963,232)(963,208)(963,208)(963,200){1}
wire w14;    //: /sn:0 {0}(719,433)(719,407)(991,407)(991,256)(974,256){1}
wire w11;    //: /sn:0 {0}(689,433)(689,371)(767,371)(767,312){1}
wire w2;    //: /sn:0 {0}(581,232)(581,170){1}
wire w15;    //: /sn:0 {0}(435,232)(435,200){1}
wire w38;    //: /sn:0 {0}(797,256)(832,256){1}
wire w43;    //: /sn:0 {0}(888,256)(918,256){1}
wire w9;    //: /sn:0 {0}(669,433)(669,371)(592,371)(592,312){1}
wire w40;    //: /sn:0 {0}(877,232)(877,200){1}
//: enddecls

  myFA g8 (.in1(w25), .in0(w2), .Cin(w23), .out(w9), .Cout(w28));   //: @(567, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  assign w30 = b[4]; //: TAP g16 @(698,194) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  myFA g3 (.in1(w1), .in0(w0), .Cin(C0), .out(w3), .Cout(w4));   //: @(304, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<0 ]
  assign w25 = b[3]; //: TAP g17 @(611,194) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  assign w16 = a[1]; //: TAP g26 @(405,164) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  //: OUT g2 (out) @(679,484) /sn:0 /R:3 /w:[ 0 ]
  assign w34 = a[5]; //: TAP g23 @(756,164) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: IN g1 (b) @(251,196) /sn:0 /w:[ 17 ]
  assign w0 = a[0]; //: TAP g24 @(318,164) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  //: IN g29 (C0) @(252,256) /sn:0 /w:[ 1 ]
  assign w20 = b[2]; //: TAP g18 @(523,194) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  myFA g10 (.in1(w35), .in0(w34), .Cin(w33), .out(w11), .Cout(w38));   //: @(742, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<0 ]
  assign w19 = a[2]; //: TAP g25 @(493,164) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  myFA g6 (.in1(w15), .in0(w16), .Cin(w4), .out(w6), .Cout(w18));   //: @(391, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  myFA g9 (.in1(w30), .in0(w17), .Cin(w28), .out(w10), .Cout(w33));   //: @(654, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<1 ]
  myFA g7 (.in1(w20), .in0(w19), .Cin(w18), .out(w8), .Cout(w23));   //: @(479, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  assign w39 = a[6]; //: TAP g22 @(847,164) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  myFA g12 (.in1(w45), .in0(w44), .Cin(w43), .out(w13), .Cout(w14));   //: @(919, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<1 ]
  assign w17 = a[4]; //: TAP g28 @(668,164) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  assign w40 = b[6]; //: TAP g14 @(877,194) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  myFA g11 (.in1(w40), .in0(w39), .Cin(w38), .out(w12), .Cout(w43));   //: @(833, 233) /sz:(54, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  assign out = {w14, w13, w12, w11, w10, w9, w8, w6, w3}; //: CONCAT g5  @(679,438) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:1
  assign w44 = a[7]; //: TAP g21 @(933,164) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  assign w15 = b[1]; //: TAP g19 @(435,194) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  assign w1 = b[0]; //: TAP g20 @(348,194) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  assign w35 = b[5]; //: TAP g15 @(786,194) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: IN g0 (a) @(250,166) /sn:0 /w:[ 17 ]
  assign w2 = a[3]; //: TAP g27 @(581,164) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  assign w45 = b[7]; //: TAP g13 @(963,194) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin myHA
module myHA(Cout, in1, out, in0);
//: interface  /sz:(48, 78) /bd:[ Ti0>in1(33/48) Ti1>in0(11/48) Bo0<out(18/48) Ro0<Cout(24/78) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(150,145)(116,145)(116,72){1}
//: {2}(118,70)(131,70){3}
//: {4}(114,70)(97,70)(97,70)(74,70){5}
input in0;    //: /sn:0 {0}(150,113)(96,113)(96,40){1}
//: {2}(98,38)(118,38)(118,38)(131,38){3}
//: {4}(94,38)(72,38){5}
output out;    //: /sn:0 {0}(185,68)(186,68)(186,68)(232,68){1}
output Cout;    //: /sn:0 {0}(206,144)(198,144)(198,144)(237,144){1}
//: enddecls

  myEXOR g4 (.in1(in1), .in0(in0), .out(out));   //: @(132, 26) /sz:(52, 55) /sn:0 /p:[ Li0>3 Li1>3 Ro0<0 ]
  //: OUT g3 (Cout) @(234,144) /sn:0 /w:[ 1 ]
  //: IN g2 (in1) @(72,70) /sn:0 /w:[ 5 ]
  //: OUT g1 (out) @(229,68) /sn:0 /w:[ 1 ]
  //: joint g6 (in0) @(96, 38) /w:[ 2 -1 4 1 ]
  //: joint g7 (in1) @(116, 70) /w:[ 2 -1 4 1 ]
  myAND g5 (.in0(in0), .in1(in1), .out(Cout));   //: @(151, 105) /sz:(54, 51) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: IN g0 (in0) @(70,38) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin REG4bit
module REG4bit(clk, out, in);
//: interface  /sz:(68, 66) /bd:[ Ti0>in[3:0](33/68) Li0>clk(45/66) Bo0<out[3:0](32/68) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] in;    //: /sn:0 {0}(#:181,238)(241,238)(241,238)(298,238){1}
//: {2}(299,238)(386,238){3}
//: {4}(387,238)(482,238){5}
//: {6}(483,238)(576,238){7}
//: {8}(577,238)(606,238){9}
output [3:0] out;    //: /sn:0 {0}(421,471)(421,448)(420,448)(#:420,443){1}
input clk;    //: /sn:0 {0}(210,268)(234,268)(234,268)(260,268){1}
//: {2}(264,268)(305,268)(305,268)(348,268){3}
//: {4}(352,268)(444,268){5}
//: {6}(448,268)(540,268)(540,312){7}
//: {8}(446,270)(446,311){9}
//: {10}(350,270)(350,312){11}
//: {12}(262,270)(262,280)(262,280)(262,311){13}
wire w6;    //: /sn:0 {0}(387,242)(387,312){1}
wire w0;    //: /sn:0 {0}(577,242)(577,312){1}
wire w3;    //: /sn:0 {0}(483,242)(483,311){1}
wire w8;    //: /sn:0 {0}(359,377)(359,408)(415,408)(415,437){1}
wire w2;    //: /sn:0 {0}(549,377)(549,422)(435,422)(435,437){1}
wire w11;    //: /sn:0 {0}(271,376)(271,422)(405,422)(405,437){1}
wire w5;    //: /sn:0 {0}(455,376)(455,408)(425,408)(425,437){1}
wire w9;    //: /sn:0 {0}(299,242)(299,250)(299,250)(299,311){1}
//: enddecls

  FFDet g4 (.clk(clk), .D(w3), .q(w5));   //: @(432, 312) /sz:(69, 63) /R:3 /sn:0 /p:[ Ti0>9 Ti1>1 Bo0<0 ]
  assign w3 = in[2]; //: TAP g8 @(483,236) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  FFDet g3 (.clk(clk), .D(w0), .q(w2));   //: @(526, 313) /sz:(69, 63) /R:3 /sn:0 /p:[ Ti0>7 Ti1>1 Bo0<0 ]
  //: IN g2 (clk) @(208,268) /sn:0 /w:[ 0 ]
  //: OUT g1 (out) @(421,468) /sn:0 /R:3 /w:[ 0 ]
  assign w9 = in[0]; //: TAP g10 @(299,236) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  FFDet g6 (.clk(clk), .D(w9), .q(w11));   //: @(248, 312) /sz:(69, 63) /R:3 /sn:0 /p:[ Ti0>13 Ti1>1 Bo0<0 ]
  assign w0 = in[3]; //: TAP g7 @(577,236) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w6 = in[1]; //: TAP g9 @(387,236) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g12 (clk) @(350, 268) /w:[ 4 -1 3 10 ]
  FFDet g5 (.clk(clk), .D(w6), .q(w8));   //: @(336, 313) /sz:(69, 63) /R:3 /sn:0 /p:[ Ti0>11 Ti1>1 Bo0<0 ]
  //: joint g11 (clk) @(446, 268) /w:[ 6 -1 5 8 ]
  assign out = {w2, w5, w8, w11}; //: CONCAT g14  @(420,442) /sn:0 /R:3 /w:[ 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  //: IN g0 (in) @(179,238) /sn:0 /w:[ 0 ]
  //: joint g13 (clk) @(262, 268) /w:[ 2 -1 1 12 ]

endmodule
//: /netlistEnd

//: /netlistBegin REG8bit
module REG8bit(out, clk, in);
//: interface  /sz:(63, 64) /bd:[ Ti0>in[7:0](30/66) Li0>clk(50/64) Ro0<out[7:0](15/64) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] in;    //: /sn:0 {0}(#:216,138)(328,138){1}
//: {2}(329,138)(371,138)(371,138)(413,138){3}
//: {4}(414,138)(497,138){5}
//: {6}(498,138)(539,138)(539,138)(579,138){7}
//: {8}(580,138)(620,138)(620,138)(659,138){9}
//: {10}(660,138)(699,138)(699,138)(738,138){11}
//: {12}(739,138)(820,138){13}
//: {14}(821,138)(859,138)(859,138)(897,138){15}
//: {16}(898,138)(919,138){17}
input clk;    //: /sn:0 {0}(222,185)(290,185){1}
//: {2}(294,185)(375,185){3}
//: {4}(379,185)(419,185)(419,185)(459,185){5}
//: {6}(463,185)(541,185){7}
//: {8}(545,185)(621,185){9}
//: {10}(625,185)(700,185){11}
//: {12}(704,185)(782,185){13}
//: {14}(786,185)(861,185)(861,213){15}
//: {16}(784,187)(784,197)(784,197)(784,213){17}
//: {18}(702,187)(702,197)(702,197)(702,213){19}
//: {20}(623,187)(623,197)(623,197)(623,213){21}
//: {22}(543,187)(543,213){23}
//: {24}(461,187)(461,197)(461,197)(461,213){25}
//: {26}(377,187)(377,213){27}
//: {28}(292,187)(292,213){29}
output [7:0] out;    //: /sn:0 {0}(589,442)(#:589,402){1}
wire w13;    //: /sn:0 {0}(564,396)(564,365)(386,365)(386,278){1}
wire w16;    //: /sn:0 {0}(574,396)(574,356)(470,356)(470,278){1}
wire w4;    //: /sn:0 {0}(594,396)(594,350)(632,350)(632,278){1}
wire w25;    //: /sn:0 {0}(604,396)(604,358)(711,358)(711,278){1}
wire w0;    //: /sn:0 {0}(624,396)(624,376)(870,376)(870,278){1}
wire w20;    //: /sn:0 {0}(660,142)(660,150)(660,150)(660,213){1}
wire w29;    //: /sn:0 {0}(898,142)(898,150)(898,150)(898,213){1}
wire w19;    //: /sn:0 {0}(584,396)(584,350)(552,350)(552,278){1}
wire w10;    //: /sn:0 {0}(554,396)(554,375)(301,375)(301,278){1}
wire w23;    //: /sn:0 {0}(739,142)(739,150)(739,150)(739,213){1}
wire w1;    //: /sn:0 {0}(614,396)(614,368)(793,368)(793,278){1}
wire w17;    //: /sn:0 {0}(580,142)(580,150)(580,150)(580,213){1}
wire w14;    //: /sn:0 {0}(498,142)(498,213){1}
wire w2;    //: /sn:0 {0}(329,142)(329,213){1}
wire w11;    //: /sn:0 {0}(414,142)(414,150)(414,150)(414,213){1}
wire w26;    //: /sn:0 {0}(821,142)(821,213){1}
//: enddecls

  FFDet g4 (.clk(clk), .D(w2), .q(w10));   //: @(278, 214) /sz:(69, 63) /R:3 /sn:0 /p:[ Ti0>29 Ti1>1 Bo0<1 ]
  FFDet g8 (.clk(clk), .D(w20), .q(w4));   //: @(609, 214) /sz:(69, 63) /sn:0 /p:[ Ti0>21 Ti1>1 Bo0<1 ]
  assign out = {w0, w1, w25, w4, w19, w16, w13, w10}; //: CONCAT g3  @(589,401) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:1
  //: joint g16 (clk) @(623, 185) /w:[ 10 -1 9 20 ]
  assign w26 = in[6]; //: TAP g26 @(821,136) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  //: joint g17 (clk) @(702, 185) /w:[ 12 -1 11 18 ]
  //: OUT g2 (out) @(589,439) /sn:0 /R:3 /w:[ 0 ]
  assign w17 = in[3]; //: TAP g23 @(580,136) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: IN g1 (clk) @(220,185) /sn:0 /w:[ 0 ]
  assign w20 = in[4]; //: TAP g24 @(660,136) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  //: joint g18 (clk) @(784, 185) /w:[ 14 -1 13 16 ]
  FFDet g10 (.clk(clk), .D(w26), .q(w1));   //: @(770, 214) /sz:(69, 63) /sn:0 /p:[ Ti0>17 Ti1>1 Bo0<1 ]
  assign w23 = in[5]; //: TAP g25 @(739,136) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  FFDet g6 (.clk(clk), .D(w14), .q(w16));   //: @(447, 214) /sz:(69, 63) /sn:0 /p:[ Ti0>25 Ti1>1 Bo0<1 ]
  FFDet g7 (.clk(clk), .D(w17), .q(w19));   //: @(529, 214) /sz:(69, 63) /sn:0 /p:[ Ti0>23 Ti1>1 Bo0<1 ]
  FFDet g9 (.clk(clk), .D(w23), .q(w25));   //: @(688, 214) /sz:(69, 63) /sn:0 /p:[ Ti0>19 Ti1>1 Bo0<1 ]
  assign w14 = in[2]; //: TAP g22 @(498,136) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g12 (clk) @(292, 185) /w:[ 2 -1 1 28 ]
  FFDet g5 (.clk(clk), .D(w11), .q(w13));   //: @(363, 214) /sz:(69, 63) /sn:0 /p:[ Ti0>27 Ti1>1 Bo0<1 ]
  FFDet g11 (.clk(clk), .D(w29), .q(w0));   //: @(847, 214) /sz:(69, 63) /sn:0 /p:[ Ti0>15 Ti1>1 Bo0<1 ]
  //: joint g14 (clk) @(461, 185) /w:[ 6 -1 5 24 ]
  assign w29 = in[7]; //: TAP g19 @(898,136) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign w11 = in[1]; //: TAP g21 @(414,136) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w2 = in[0]; //: TAP g20 @(329,136) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: IN g0 (in) @(214,138) /sn:0 /w:[ 0 ]
  //: joint g15 (clk) @(543, 185) /w:[ 8 -1 7 22 ]
  //: joint g13 (clk) @(377, 185) /w:[ 4 -1 3 26 ]

endmodule
//: /netlistEnd

